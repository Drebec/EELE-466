library IEEE;
use IEEE.std_logic_1164.all;

entity four_bit_cla_adder is
  port( A, B 	: in std_logic_vector(3 downto 0);
	Cin  	: in std_logic;
	S 	: out std_logic_vector(3 downto 0);
	Cout 	: out std_logic);
end entity;

architecture four_bit_cla_adder_arch of four_bit_cla_adder is

  signal P, G, C : std_logic_vector(3 downto 0);

  begin

  P(0) <= A(0) xor B(0);
  P(1) <= A(1) xor B(1);
  P(2) <= A(2) xor B(2);
  P(3) <= A(3) xor B(3);

  G(0) <= A(0) and B(0);
  G(1) <= A(1) and B(1);
  G(2) <= A(2) and B(2);
  G(3) <= A(3) and B(3);

  C(0) <= Cin;
  C(1) <= G(0) or (P(0) and C(0));
  C(2) <= G(1) or (P(1) and C(1));
  C(3) <= G(2) or (P(2) and C(2));
  Cout <= G(3) or (P(3) and C(3));

  S(0) <= P(0) xor C(0);
  S(1) <= P(1) xor C(1);
  S(2) <= P(2) xor C(2);
  S(3) <= P(3) xor C(3);

end architecture;
